module top_tb;
    import uvm_pkg::*;
    initial begin
        #1ns;
        `uvm_info("soc_top_tb", "******************************************************************************", UVM_NONE)
        `uvm_info("soc_top_tb", "**************************in soc_top_tb for default **************************", UVM_NONE)
        `uvm_info("soc_top_tb", "******************************************************************************", UVM_NONE)
    end
endmodule
